module rom(address,data);
	input [8:0] address; //needs to be changed
	output [60:0] data;	//needs to be changed
	reg [60:0] array[511:0];	//needs to be changed
	always @*
		begin

			/*** NOP ***/
			array[0] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION
			/*** 25_NOP ***/
			array[320] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000001_000_000; // cycle until i say
			array[321] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000010_000_000; // cycle until i say
			array[322] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000011_000_000; // cycle until i say
			array[323] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000100_000_000; // cycle until i say
			array[324] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000101_000_000; // cycle until i say
			array[325] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000110_000_000; // cycle until i say
			array[326] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101000111_000_000; // cycle until i say
			array[327] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001000_000_000; // cycle until i say
			array[328] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001001_000_000; // cycle until i say
			array[329] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001010_000_000; // cycle until i say
			array[330] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001011_000_000; // cycle until i say
			array[331] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001100_000_000; // cycle until i say
			array[332] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001101_000_000; // cycle until i say
			array[333] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001110_000_000; // cycle until i say
			array[334] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101001111_000_000; // cycle until i say
			array[335] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010000_000_000; // cycle until i say
			array[336] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010001_000_000; // cycle until i say
			array[337] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010010_000_000; // cycle until i say
			array[338] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010011_000_000; // cycle until i say
			array[339] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010100_000_000; // cycle until i say
			array[340] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010101_000_000; // cycle until i say
			array[341] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010110_000_000; // cycle until i say
			array[342] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_101010111_000_000; // cycle until i say
			array[343] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_001000000000_0_0_100001100_000_000; // cycle until i say
			//array[344] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1101_0000_001000000000_0_0_100001100_000_000; // cycle until i say
			/** BIPUSH **/
			array[16] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000010000000_1_0_000010001_000_000; // ORS <- MDR_rd >> 8
			array[17] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_100000001000_0_0_000010010_000_000; // MAR <- SP <- SP + 4
			array[18] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0001_0000_001000000000_0_0_000010100_000_000; // MDR_wr <- ORS
			array[20] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000011101_101_000; // START, WRITE
			array[29] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** LDC_W **/ 
			array[19] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000010000001_1_0_000001111_000_000; // EXR <- ORS <- MDR_RD >> 8, PC++
			array[15] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000001000000_1_0_000000001_000_000; // ORU <- EXR >> 8, PC++
			array[1] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_0001_0000_000000000010_0_0_000000010_000_000; // TMR <- ORS << 8
			array[2] = 61'b0_0_0_000_000_0_0_0_0_011100_0010_0_0111_0010_000000000010_0_0_000000011_000_000; // TMR <- TMR OR ORU << 2
			array[3] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0111_0110_100000000000_0_0_000000100_000_000; // MAR <- CPP + TMR
			array[4] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_000000001000_0_0_000000101_110_000; // START, READ, SP <- SP + 4
			array[5] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_110000000000_0_0_000000110_000_000; // MDR_RD <- MEM_READ, MAR <- SP
			array[6] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_000000111_000_000; // MDR_WR <- MDR_RD
			array[7] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000001000_101_000; // START, WRITE
			array[8] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** ILOAD **/
			array[21] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000001000000_1_0_000010110_000_000; // ORU <- MDR_rd >> 8, PC++
			array[22] = 61'b0_0_0_000_000_0_0_0_0_011000_0010_0_0010_0000_000001000000_0_0_000010111_000_000; // ORU <- ORU << 2
			array[23] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0100_0010_100000000000_0_0_000011000_000_000; // MAR <- LV + ORU
			array[24] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_000000001000_0_0_000011001_110_000; // START, RWN, SP <- SP + 4
			array[25] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_110000000000_0_0_000011010_000_000; // MDR_rd <- MEM_read, MAR <- SP
			array[26] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_000011011_000_000; // MDR_wr <- MDR_rd
			array[27] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000011100_101_000; // START, WRITE
			array[28] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** ISTORE **/
			array[54] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000001000000_0_0_000110111_000_000; // ORU <- MDR >> 8
			array[55] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_000111000_000_000; // MAR <- SP
			array[56] = 61'b0_0_0_000_000_0_0_0_0_011000_0010_0_0010_0000_000000000010_0_0_000111001_110_000; // START, RWN, TMR <- ORU << 2
			array[57] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0100_0111_110000000000_0_0_000111010_000_000; // MDR_rd <- MEM_read, MAR <- LV + TMR
			array[58] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_000111011_000_000; // MDR_wr <- MDR_rd
			array[59] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_1_0_000111100_101_000; // START, SP <- SP - 4, PC++
			array[60] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** POP **/
			array[87] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_100000000_000_000; // SP <- SP - 4, GOTO CYCLE_DECISION

			/** DUP **/
			array[89] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_001011010_000_000; // MAR <- SP
			array[90] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_000000001000_0_0_001011011_110_000; // START, READ, SP <- SP + 4
			array[91] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_110000000000_0_0_001011100_000_000; // MDR_rd <- MEM_READ, MAR <- SP
			array[92] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_001011101_000_000; // MDR_wr <- MDR_rd
			array[93] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001011110_101_000; // START, WRITE
			array[94] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** SWAP **/
			array[95] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_001000000_000_000; // MAR <- SP
			array[64] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001000001_110_000; // START, READ
			array[65] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_110000000000_0_0_001000010_000_000; // MDR_rd <- MEM_read, MAR <- SP - 4
			array[66] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000010_0_0_001000011_110_000; // START, READ, TMR <- MDR_rd
			array[67] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0111_0000_011000000000_0_0_001000100_000_000; // MDR_rd <- MEM_read, MDR_wr <- TMR
			array[68] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001000101_101_000; // START, WRITE
			array[69] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_001000110_000_000; // MDR_wr <- MDR_rd
			array[70] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_001000111_000_000; // MAR <- SP
			array[71] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001001000_101_000; // START, WRITE
			array[72] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** IADD **/
			array[96] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_001100001_000_000; // MAR <- SP
			array[97] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001100010_110_000; // START, READ
			array[98] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_110000000000_0_0_001100011_000_000; // MDR_rd <- MEM_read, MAR <- SP - 4
			array[99] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_001100101_110_000; // START, READ, SP <- SP - 4
			array[101] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_010000000010_0_0_001100110_000_000; // MDR_rd <- MEM_read, TMR <- MDR_rd
			array[102] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0000_0111_001000000000_0_0_001100111_000_000; // MDR_wr <- MDR_rd + TMR
			array[103] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001101000_101_000; // START, WRITE
			array[104] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** ISUB **/
			array[100] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_001101001_000_000; // MAR <- SP
			array[105] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001101010_110_000; // START, READ
			array[106] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_110000000000_0_0_001101011_000_000; // MDR_rd <- MEM_read, MAR <- SP - 4
			array[107] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_001101100_110_000; // START, READ, SP <- SP - 4
			array[108] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_010000000010_0_0_001101101_000_000; // MDR_rd <- MEM_read, TMR <- MDR_rd
			array[109] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_0000_0111_001000000000_0_0_001101110_000_000; // MDR_wr <- MDR_rd - TMR
			array[110] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001110000_101_000; // START, WRITE
			array[112] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** IAND **/
			array[126] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_001110001_000_000; // MAR <- SP
			array[113] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001110010_110_000; // START, READ
			array[114] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_110000000000_0_0_001110011_000_000; // MDR_rd <- MEM_read, MAR <- SP - 4
			array[115] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_001110100_110_000; // START, READ, SP <- SP - 4
			array[116] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_010000000010_0_0_001110101_000_000; // MDR_rd <- MEM_read, TMR <- MDR_rd
			array[117] = 61'b0_0_0_000_000_0_0_0_0_001100_0000_0_0000_0111_001000000000_0_0_001110110_000_000; // MDR_wr <- MDR_rd AND TMR
			array[118] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001110111_101_000; // START, WRITE
			array[119] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** IOR **/
			array[128] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_010000001_000_000; // MAR <- SP
			array[129] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010000010_110_000; // START, READ
			array[130] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_110000000000_0_0_010000011_000_000; // MDR_rd <- MEM_read, MAR <- SP - 4
			array[131] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_001111000_110_000; // START, READ, SP <- SP - 4
			array[120] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_010000000010_0_0_001111001_000_000; // MDR_rd <- MEM_read, TMR <- MDR_rd
			array[121] = 61'b0_0_0_000_000_0_0_0_0_011100_0000_0_0000_0111_001000000000_0_0_001111010_000_000; // MDR_wr <- MDR_rd OR TMR
			array[122] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001111011_101_000; // START, WRITE
			array[123] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** IINC **/
			array[132] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000001000010_1_0_010000101_000_000; // ORU <- TMR <- MDR_rd >> 8
			array[133] = 61'b0_0_0_000_000_0_0_0_0_011000_0010_0_0010_0000_000001000000_1_0_010000110_000_000; // ORU <- ORU << 2
			array[134] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0010_0100_100000000000_0_0_010000111_000_000; // MAR <- ORU + LV
			array[135] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0111_0000_000010000000_0_0_010001000_110_000; // START, READ, ORS <- TMR >> 8
			array[136] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_010001001_000_000; // MDR_rd <- MEM_read
			array[137] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0000_0001_001000000000_0_0_010001010_000_000; // MDR_wr <- MDR_rd + ORS
			array[138] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010001011_101_000; // START, WRITE
			array[139] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** IFEQ **/
			array[153] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_010010111_000_000; // MAR <- SP
			array[151] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_010011010_000_000; // SP <- SP - 4
			array[154] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000001_0_0_010011100_110_000; // START, READ, EXR <- MDR_rd
			array[156] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_010011101_000_000; // MDR_rd <- MEM_read
			array[157] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000010_0_0_010011110_000_001; // TMR <- MDR_rd
			array[158] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_1_0_010011000_000_000; // PC++
			array[152] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_1_0_100000000_000_000; // PC++, GOTO CYCLE_DECISION
			array[414] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010101000_000_000; // GOTO GOTO

			/** IFLT **/
			array[155] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_011010000_000_000; // MAR <- SP
			array[208] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_011010001_000_000; // SP <- SP - 4
			array[209] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000001_0_0_011010010_110_000; // START, READ, EXR <- MDR_rd
			array[210] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_011010011_000_000; // MDR_rd <- MEM_read
			array[211] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000010_0_0_011010100_000_010; // TMR <- MDR_rd
			array[212] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_1_0_011010101_000_000; // PC++
			array[213] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_1_0_011010110_000_000; // PC++
			array[468] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010101000_000_000; // GOTO GOTO

			/** IF_ICMPEQ **/
			array[159] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_011011111_000_000; // MAR <- SP
			array[223] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_011100000_000_000; // SP <- SP - 4
			array[224] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000001_0_0_011100001_110_000; // START, READ, EXR <- MDR_rd
			array[225] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_110000000000_0_0_011100010_000_000; // MDR_rd <- MEM_read, MAR <- SP
			array[226] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000010_0_0_011100011_110_000; // START, READ, TMR <- MDR_rd
			array[227] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_011011110_000_000; // MDR_rd <- MEM_read
			array[222] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_011100100_000_000; // SP <- SP - 4
			array[228] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_0000_0111_000000000010_0_0_011100101_000_001; // TMR <- TMR - MDR_rd
			array[229] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_1_0_011100110_000_000; // PC++
			array[230] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_1_0_100000000_000_000; // PC++, GOTO CYCLE_DECISION
			array[485] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010101000_000_000; // GOTO GOTO 

			/** GOTO **/
			array[167] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000001_0_0_010101000_000_000; // EXR <- MDR_rd

			array[168] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000010000001_0_0_010101001_000_000; // ORS <- EXR >> 8, EXR <- EXR >> 8
			array[169] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000001000001_0_0_010101010_000_000; // ORU <- EXR >> 8
			array[170] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_0001_0000_000000000010_0_0_010101011_000_000; // TMR <- ORS << 8
			array[171] = 61'b0_0_0_000_000_0_0_0_0_011100_0000_0_0111_0010_000000000010_0_0_010101101_000_000; // TMR <- ORU OR TMR

			array[173] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0011_0111_000000100000_0_0_010101110_000_000; // PC <- PC + TMR
			array[174] = 61'b0_0_0_000_000_0_0_0_0_110110_0000_0_0000_0011_000000100000_0_0_100000000_000_000; // PC <- PC - 1

			/** INVOKE **/
			array[182] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000000001_1_0_010110111_000_000; // EXR <- MDR_rd
			array[183] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000010000001_1_0_010111000_000_000; // EXR <- ORS <- EXR >> 8
			array[184] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000001000000_0_0_010111001_000_000; // ORU <- EXR >> 8
			array[185] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_0001_0000_000000000010_0_0_010111010_000_000; // TMR <- ORS << 8
			array[186] = 61'b0_0_0_000_000_0_0_0_0_011100_0010_0_0111_0010_000000000010_0_0_010111011_000_000; // TMR <- (ORU OR TMR) << 2
			array[187] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0111_0110_100000000000_0_0_010111100_000_000; // MAR <- CPP + TMR

			array[188] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010111101_110_000; // START, READ
			array[189] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_010111110_000_000; // MDR_rd <- MEM_read
 			array[190] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_100000000100_0_0_010111111_000_000; // MAR <- CPP <- MDR_rd
 			array[191] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_011111111_110_000; // START, READ
 			array[255] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_011000000_000_000; // MDR_rd <- MEM_read
 			array[192] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_0000_0000_000000000001_0_0_011000001_000_000; // EXR <- MDR_rd << 8
 			array[193] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_1000_0000_000000000001_0_0_011000010_000_000; // EXR <- EXR << 8
 			array[194] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000000000001_0_0_011000011_000_000; // EXR <- EXR >> 8
 			array[195] = 61'b0_0_0_000_000_0_0_0_0_011000_0110_1_1000_0000_000000000001_0_0_011000110_000_000; // EXR <- EXR >> 6
 			array[198] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1000_0101_000000000001_0_0_011000111_000_000; // EXR <- SP - EXR
 			array[199] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000000000010_0_0_011001000_000_000; // TMR <- MDR_rd >> 8
 			array[200] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0111_0000_000000000010_0_0_011001001_000_000; // TMR <- TMR >> 8
 			array[201] = 61'b0_0_0_000_000_0_0_0_0_011000_0010_0_0111_0000_000000000010_0_0_011001010_000_000; // TMR <- TMR << 2
 			array[202] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1000_0000_100000000000_0_0_011001011_000_000; // MAR <- EXR
 			array[203] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0111_0101_000000000010_0_0_011001100_000_000; // TMR <- SP + TMR
 			array[204] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0111_001000000010_0_0_011001101_000_000; // MDR_wr <- TMR <- TMR + CONST4
 			array[205] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_011001110_101_000; // START, WRITE
 			array[206] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0111_0000_100000001000_0_0_011001111_000_000; // MAR <- SP <- TMR
 			array[207] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0011_0000_001000000000_0_0_011110000_000_000; // MDR_wr <- PC
 			array[240] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0101_1001_000000001000_0_0_011110001_101_000; // START, WRITE, SP <- SP + CONST4
 			array[241] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_011110010_000_000; // MAR <- SP
 			array[242] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0100_0000_001000000000_0_0_011110011_000_000; // MDR_wr <- LV
 			array[243] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_011110100_101_000; // START, WRITE
 			array[244] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1000_0000_000000010000_0_0_011110101_000_000; // LV <- EXR
 			array[245] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0110_1001_000000100000_0_0_011110110_000_000; // PC <- CPP + CONST4
 			array[246] = 61'b0_0_0_000_000_0_0_0_0_110001_0110_0_0000_0000_000000000100_0_0_100000000_000_000; // CPP <- 1 << 6, GOTO CYCLE_DECISION

 			/** IRETURN **/ 
 			array[172] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0100_0000_100000001000_0_0_010101101_000_000; // MAR <- SP <- LV
 			array[173] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010101110_110_000; // START, READ
 			array[174] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_010101111_000_000; // MDR_rd <- MEM_read
 			array[175] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_100000000010_0_0_010110000_000_000; // MAR <- TMR <- MDR_rd
 			array[176] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010110001_110_000; // START, READ
 			array[177] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_010110010_000_000; // MDR_rd <- MEM_read
 			array[178] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000100000_0_0_010110011_000_000; // PC <- MDR_rd
 			array[179] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0111_1001_100000000010_0_0_010110100_000_000; // MAR <- TMR + CONST4
 			array[180] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_010110101_110_000; // START, READ
 			array[181] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_011110111_000_000; // MDR_rd <- MEM_read
 			array[247] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000000010000_0_0_011111000_000_000; // LV <- MDR_rd
 			array[248] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0111_100000000000_0_0_011111001_000_000; // MAR <- TMR + CONST4
 			array[249] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_011111010_110_000; // START, READ
 			array[250] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_011111011_000_000; // MDR_rd <- MEM_read
 			array[251] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_011111100_000_000; // MDR_wr <- MDR_rd
 			array[252] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_011111101_000_000; // MAR <- SP
 			array[253] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_011111110_101_000; // START, READ
 			array[254] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** WIDE **/
			array[196] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000100000001_1_0_011000101_000_000; // IR <- EXR <- MDR_rd >> 8, PC++
			array[197] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_1_000000000_000_100; // GOTO WIDE_OPCODE

			/** FETCH **/
			array[511] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0011_0000_100000000000_1_0_100000001_000_000; // MAR <- PC, PC++
			array[257] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000010_110_000; // START, READ
			array[258] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_100000011_000_000; // MDR_rd <- MEM_read
			array[259] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_000100000000_0_0_100000100_000_000; // IR <- OPCODE
			array[260] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000000000_000_100; // GOTO OPCODE

			/** WIDE_ISTORE **/
			array[310] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000000000001_1_0_100110111_000_000; // EXR <- EXR >> 8, PC++
			array[311] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000001000000_1_0_100111000_000_000; // ORU <- EXR << 8, PC++
			array[312] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_1000_0000_000000000010_0_0_100111001_000_000; // TMR <- EXR >> 8
			array[313] = 61'b0_0_0_000_000_0_0_0_0_011100_0010_0_0111_0010_000000000010_0_0_100111010_000_000; // TMR <- TMR OR ORU
			array[314] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_100111011_000_000; // MAR <- SP
			array[315] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100111100_110_000; // START, READ
			array[316] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0111_0100_110000000000_0_0_100111101_000_000; // MDR_rd <- MEM_read, MAR <- TMR + LV
			array[317] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_100111110_000_000; // MDR_wr <- MDR_rd
			array[318] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_100111111_101_000; // START, WRITE, SP <- SP - 4
			array[319] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION

			/** WIDE_ILOAD **/
			array[277] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000000000001_1_0_100010110_000_000; // EXR <- EXR >> 8
			array[278] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_1000_0000_000001000000_1_0_100010111_000_000; // ORU <- EXR >> 8
			array[279] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_0_1000_0000_000000000010_0_0_100011000_000_000; // TMR <- EXR << 8
			array[280] = 61'b0_0_0_000_000_0_0_0_0_011100_0010_0_0111_0010_000000000010_0_0_100011001_000_000; // TMR <- (TMR OR ORU) << 2
			array[281] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_0100_0111_100000000000_0_0_100011010_000_000; // MAR <- LV + TMR 
			array[282] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_000000001000_0_0_100011011_110_000; // START, READ, SP <- SP + CONST4
			array[283] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_110000000000_0_0_100011100_000_000; // MDR_rd <- MEM_read, MAR <- SP
			array[284] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_001000000000_0_0_100011101_000_000; // MDR_wr <- MDR_rd
			array[285] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100011110_101_000; // START, WRITE
			array[286] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION
			
			/** INPUT **/
			array[9] = 61'b0_0_0_000_100_0_0_0_1_000000_0000_0_1010_0000_000011000000_0_0_000001010_000_000; // ORS <- ORU <- IO_INPUT
			array[10] = 61'b0_0_0_000_100_0_0_0_1_000000_0000_0_1010_0000_001000000000_0_0_100000000_000_000; // MDR_wr <- IO_INPUT
			array[11] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_100000001000_0_0_000011111_000_000; // MAR <- SP <- SP + 4
			array[12] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000100111_101_000; // START, WRITE
			array[13] = 61'b0_0_0_000_100_1_1_0_1_000000_0000_0_1010_0000_000011000000_0_0_100000000_000_000; // TOGGLE IE, GOTO CYCLE_DECISION
			
			/** CYCLE_DECISION **/
			array[256] = 61'b0_0_1_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_111111111_000_000; // If interrupt GOTO INTERRUPT_CHECK Else GOTO FETCH
			
			/** INTERRUPT_CHECK **/
			array[125] = 61'b0_0_0_000_010_0_0_0_0_011000_1000_1_1011_1010_000010000000_1_0_001111111_000_000; // if interrupt_level - PIL < 0 SKIP NEXT LINE
			array[127] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_111111111_000_000; // GOTO FETCH
			array[383] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000001110_000_000; // GOTO INTERRUPT
			
			/** INTERRUPT **/
			array[30] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_100000001000_0_0_000011111_000_000; // MAR <- SP <- SP + 4
			array[31] = 61'b0_0_0_000_001_0_0_0_0_011000_0000_0_1010_0000_001000000000_0_0_000100000_000_000; // MDR_wr <- PSR
			array[32] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000100001_101_000; // START, WRITE
			
			array[33] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_100000001000_0_0_000100010_000_000; // MAR <- SP <- SP + 4
			array[34] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0011_0000_001000000000_0_0_000100011_000_000; // MDR_wr <- PC
			array[35] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000100100_101_000; // START, WRITE
			
			array[36] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_100000001000_0_0_000100101_000_000; // MAR <- SP <- SP + 4
			array[37] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1100_0000_001000000000_0_0_000100110_000_000; // MDR_wr <- FRAME
			array[38] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000100111_101_000; // START, WRITE
			
			array[39] = 61'b0_0_0_000_000_0_0_0_0_111100_0000_0_1001_0101_100000001000_0_0_000101000_000_000; // MAR <- SP <- SP + 4
			array[40] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0100_0000_001000000000_0_0_000101001_000_000; // MDR_wr <- LV
			array[41] = 61'b1_0_0_000_000_1_1_0_0_000000_0000_0_0000_0000_000000000000_0_0_000101010_101_000; // START, WRITE, IE <- 0, FRAME <- SP
			
			array[42] = 61'b1_0_0_000_000_0_0_0_1_011000_0000_0_1001_0000_000000000000_0_0_000101011_000_000; // FRAME <- SP
			array[43] = 61'b0_0_0_000_011_1_1_1_1_011000_0000_0_1010_0000_100000000000_0_0_000101100_101_000; // LOAD PIL, MAR <- TRAPBASE
			array[44] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_000101101_110_000; // START, READ
			array[45] = 61'b0_0_0_000_000_0_0_0_0_011100_0000_0_0000_0000_000000100000_0_0_100000000_000_000; // PC <- MDR_RD, GOTO CYCLE_DECISION
			
			/** INT_RET **/
			array[73] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1100_0000_100000001000_0_0_001001010_000_000; // MAR <- SP <- FRAME
 			array[74] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001001011_110_000; // START, READ
 			array[75] = 61'b1_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000000000_0_0_001001100_000_000; // FRAME <- MEM_read
 			
 			array[76] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1001_0101_100000001000_0_0_001001101_000_000; // MAR <- SP <- SP - 4
 			array[77] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001001110_110_000; // START, READ
 			array[78] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000010000_0_0_001001111_000_000; // LV <- MEM_read
 			
 			array[79] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1001_0101_100000001000_0_0_001010000_000_000; // MAR <- SP <- SP - 4
 			array[80] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001010001_110_000; // START, READ
 			array[81] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_010000100000_0_0_001010010_000_000; // PC <- MEM_read
 			
 			array[82] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_1001_0101_100000001000_0_0_001010011_000_000; // MAR <- SP <- SP - 4
 			array[83] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_001010100_110_000; // START, READ
 			array[84] = 61'b0_1_0_000_000_0_0_1_0_000000_0000_0_0000_0000_010000000000_0_0_001010101_000_000; // PSR <- MEM_read
 			
 			array[85] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_100000000_000_000; // SP <- SP - 4
			/** floating point mult **/
			array[261] = 61'b0_0_0_000_000_0_0_0_0_011000_1000_1_0000_0000_000010000000_1_0_100000110_000_000; // ORS <- MDR_rd >> 8
			array[262] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0101_0000_100000000000_0_0_100000111_000_000; // MAR <- SP
			array[263] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100001000_110_000; // START, READ
			array[264] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_110000000000_0_0_100001001_000_000; // MDR_rd <- MEM_read, MAR <- SP - 4
			array[265] = 61'b0_0_0_000_000_0_0_0_0_111111_0000_0_1001_0101_000000001000_0_0_100001010_110_000; // START, READ, SP <- SP - 4
			array[266] = 61'b0_0_0_000_000_0_0_0_0_011000_0000_0_0000_0000_010000000010_0_0_100001011_000_000; // MDR_rd <- MEM_read, TMR <- MDR_rd
			array[267] = 61'b0_0_0_000_000_0_0_0_0_100000_0000_0_0000_0111_000000000000_0_0_101000000_000_000; // MDR_rd mult TMR
			array[268] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100001101_101_000; // START, WRITE
			array[269] = 61'b0_0_0_000_000_0_0_0_0_000000_0000_0_0000_0000_000000000000_0_0_100000000_000_000; // GOTO CYCLE_DECISION
			
		end
	assign data = array[address];
endmodule
