jjSub_inst : jjSub PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
