IR_inst : IR PORT MAP (
		clock	 => clock_sig,
		cnt_en	 => cnt_en_sig,
		data	 => data_sig,
		sclr	 => sclr_sig,
		sload	 => sload_sig,
		sset	 => sset_sig,
		q	 => q_sig
	);
