INIT_CPP_inst : INIT_CPP PORT MAP (
		result	 => result_sig
	);
