finalAdder_inst : finalAdder PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
