SpecialMantissCorrection_inst : SpecialMantissCorrection PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
