CONST4_inst : CONST4 PORT MAP (
		result	 => result_sig
	);
