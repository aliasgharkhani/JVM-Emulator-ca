CONST24_inst : CONST24 PORT MAP (
		result	 => result_sig
	);
