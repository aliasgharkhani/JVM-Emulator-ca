subtracter_inst : subtracter PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
