SHRA_inst : SHRA PORT MAP (
		data	 => data_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
