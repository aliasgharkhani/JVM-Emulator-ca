INIT_LV_inst : INIT_LV PORT MAP (
		result	 => result_sig
	);
