negativer_inst : negativer PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
