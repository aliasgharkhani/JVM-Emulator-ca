newModule_inst : newModule PORT MAP (
		dataa	 => dataa_sig,
		result	 => result_sig
	);
