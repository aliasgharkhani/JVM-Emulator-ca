negativer26bit_inst : negativer26bit PORT MAP (
		datab	 => datab_sig,
		result	 => result_sig
	);
