ALU_SHIFTER_inst : ALU_SHIFTER PORT MAP (
		data	 => data_sig,
		direction	 => direction_sig,
		distance	 => distance_sig,
		result	 => result_sig
	);
