adder_inst : adder PORT MAP (
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		overflow	 => overflow_sig,
		result	 => result_sig
	);
