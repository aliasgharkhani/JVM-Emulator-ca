INIT_SP_inst : INIT_SP PORT MAP (
		result	 => result_sig
	);
